///////////////////////
/// PACKAGE: SA_PKG ///
///////////////////////
package sa_pkg;

endpackage

////////////////////////
/// INTERFACE: PE_IF ///
////////////////////////
// interface pe_if
// #(
//     parameter ADD_DATAWIDTH,
//     parameter MUL_DATAWIDTH
// )();
//
// endinterface


import sa_pkg::*;

module sa_control
#(
    parameter ADD_DATAWIDTH,
    parameter MUL_DATAWIDTH,
    parameter NUM_ROWS,
    parameter NUM_COLS
) (
    ports
);
    
endmodule